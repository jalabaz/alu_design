library verilog;
use verilog.vl_types.all;
entity aluMain_vlg_vec_tst is
end aluMain_vlg_vec_tst;
