library verilog;
use verilog.vl_types.all;
entity ALU_DESIGN_vlg_vec_tst is
end ALU_DESIGN_vlg_vec_tst;
